module helloworld;
    initial
    begin 
    $display("Hello World!");
    $finish;
    end
endmodule
